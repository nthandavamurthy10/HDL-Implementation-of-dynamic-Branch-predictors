library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;


entity tb_onebitpred is
end tb_onebitpred;


architecture test of tb_onebitpred is 
signal branch_addr: bit;
signal branch_pred:std_logic;
signal miss_prednum:integer;

component one_bitpredictor is
port( branch_address:in bit;
      current_prediction:in std_logic;
      miss_prediction:out integer);
end component;
begin
dut: one_bitpredictor port map (branch_address => branch_addr,current_prediction => branch_pred,miss_prediction=>miss_prednum);
stimulus: process
begin
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '0';
wait for 10 ns;

wait;

end process stimulus;
end;