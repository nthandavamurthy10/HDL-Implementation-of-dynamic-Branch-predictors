library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_bit.all;
use IEEE.STD_LOGIC_ARITH.ALL;
use ieee.std_logic_unsigned.all;

entity tb_twobitpred is
end tb_twobitpred;

architecture test of tb_twobitpred is 
signal branch_addr: bit;
signal branch_pred:std_logic;
signal miss_prednum:integer:=0;

component twobit_predictor
port( b_address:in bit;
      branch_prediction:in std_logic;
      miss_prediction:out integer);
end component;
begin
dut: twobit_predictor port map (b_address => branch_addr,branch_prediction => branch_pred,miss_prediction=>miss_prednum);
stimulus: process
begin

branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '1';
wait for 10 ns;
branch_addr <= '1';
branch_pred <= '0';
wait for 10 ns;
branch_addr <= '0';
branch_pred <= '0';
wait;

end process stimulus;
end;